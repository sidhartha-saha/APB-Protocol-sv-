library verilog;
use verilog.vl_types.all;
entity apb_pkg_sv_unit is
end apb_pkg_sv_unit;
