library verilog;
use verilog.vl_types.all;
entity apb_test_sv_unit is
end apb_test_sv_unit;
