library verilog;
use verilog.vl_types.all;
entity apb_interface is
end apb_interface;
