library verilog;
use verilog.vl_types.all;
entity tb_top_sv_unit is
end tb_top_sv_unit;
