class apb_packet;
   logic [7:0] addr;
   logic [31:0] data;


endclass
